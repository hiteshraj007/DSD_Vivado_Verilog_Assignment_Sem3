`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 19.11.2025 17:30:32
// Design Name: 
// Module Name: counter_design
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module counter_design(
    input clk,
    input reset,
    input up_down,            
    output reg [3:0] count
    );
    always @(posedge clk or posedge reset) begin
    if (reset)
        count <= 0;
    else if (up_down)
        count <= count + 1;
    else
        count <= count - 1;
end
endmodule
